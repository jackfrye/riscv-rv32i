module alu
#(
  parameter integer WIDTH = 32
)
(
  input              clk        ,
  input              rst        ,
  input  [WIDTH-1:0] a          ,
  input  [WIDTH-1:0] b          ,
  input  [2:0]       alu_control,
  output [WIDTH-1:0] out
);
// STUB


endmodule